module decode (

    input logic clk;
    input logic 

);


endmodule 